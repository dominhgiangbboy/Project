library ieee;
use ieee.std_logic_1164.all;
-------------------------------------------------------
entity demux_1to32_1 is
	port(
		clk : in std_logic;
		A : in std_logic;
		sel : in std_logic_vector(4 downto 0);
		en : in std_logic := '0';
		B : out std_logic_vector(31 downto 0)
		);
end demux_1to32_1;
--------------------------------------------------------

architecture arch of demux_1to32_1 is

begin
	process(clk)
	begin
	if(en = '1') and rising_edge(clk)then
		if    sel = "11111" then B <= A & "0000000000000000000000000000000";--32
		elsif sel = "11110" then B <= '0' & A &"000000000000000000000000000000";--31
		elsif sel = "11101" then B <= "00" & A &"00000000000000000000000000000";--30
		elsif sel = "11100" then B <= "000" & A &"0000000000000000000000000000";--29
		elsif sel = "11011" then B <= "0000" & A &"000000000000000000000000000";--28
		elsif sel = "11010" then B <= "00000" & A &"00000000000000000000000000";--27
		elsif sel = "11001" then B <= "000000" & A &"0000000000000000000000000";--26
		elsif sel = "11000" then B <= "0000000" & A &"000000000000000000000000";--25
		elsif sel = "10111" then B <= "00000000" & A &"00000000000000000000000";--24
		elsif sel = "10110" then B <= "000000000" & A &"0000000000000000000000";--23
		elsif sel = "10101" then B <= "0000000000" & A &"000000000000000000000";--22
		elsif sel = "10100" then B <= "00000000000" & A &"00000000000000000000";--21
		elsif sel = "10011" then B <= "000000000000" & A &"0000000000000000000";--20
		elsif sel = "10010" then B <= "0000000000000" & A &"000000000000000000";--19
		elsif sel = "10001" then B <= "00000000000000" & A &"00000000000000000";--18
		elsif sel = "10000" then B <= "000000000000000" & A &"0000000000000000";--17
		elsif sel = "01111" then B <= "0000000000000000" & A &"000000000000000";--16
		elsif sel = "01110" then B <= "00000000000000000" & A &"00000000000000";--15
		elsif sel = "01101" then B <= "000000000000000000" & A &"0000000000000";--14
		elsif sel = "01100" then B <= "0000000000000000000" & A &"000000000000";--13
		elsif sel = "01011" then B <= "00000000000000000000" & A &"00000000000";--12
		elsif sel = "01010" then B <= "000000000000000000000" & A &"0000000000";--11
		elsif sel = "01001" then B <= "0000000000000000000000" & A &"000000000";--10
		elsif sel = "01000" then B <= "00000000000000000000000" & A &"00000000";--9
		elsif sel = "00111" then B <= "000000000000000000000000" & A &"0000000";--8
		elsif sel = "00110" then B <= "0000000000000000000000000" & A &"000000";--7
		elsif sel = "00101" then B <= "00000000000000000000000000" & A &"00000";--6
		elsif sel = "00100" then B <= "000000000000000000000000000" & A &"0000";--5
		elsif sel = "00011" then B <= "0000000000000000000000000000" & A &"000";--4
		elsif sel = "00010" then B <= "00000000000000000000000000000" & A &"00";--3
		elsif sel = "00001" then B <= "000000000000000000000000000000" & A &"0";--2
		elsif sel = "00000" then B <= "0000000000000000000000000000000" & A;--1
		end if;	
	end if;
	end process;
	
end arch;